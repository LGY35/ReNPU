module vbrain_recuc #(
    localparam DATA_FIFO_DEPTH      = 64 ,
    localparam DATA_FIFO_CNT_WID    = 6+1,
    localparam ADDR_FIFO_DEPTH      = 32 ,
    localparam ADDR_FIFO_CNT_WID    = 5+1,

    localparam D_AXI_DATA_WID       = 256,
    localparam D_AXI_ADDR_WID       = 32 ,
    localparam D_AXI_IDW            = 4  ,
    localparam D_AXI_LENW           = 4  ,
    localparam D_AXI_LOCKW          = 1  ,
    localparam D_AXI_STRBW          = 32 ,

    localparam AXI_DW               = 128,
    localparam AXI_AW               = 32,
    localparam STRB_WIDTH           = (AXI_DW/8),
    localparam ID_WIDTH             = 8,
    localparam AXI_LENW             = 4,
    localparam AXI_LOCKW            = 1,
    localparam I_FLIT_WIDTH         = 32
)
(

    input                                   clk,
    input                                   rst_n,

    //data
    output                             d_arvalid_0,
    output  [D_AXI_IDW-1:0]            d_arid_0   ,
    output  [D_AXI_ADDR_WID-1:0]       d_araddr_0 ,
    output  [D_AXI_LENW-1:0]           d_arlen_0  ,
    output  [2:0]                      d_arsize_0 ,
    output  [1:0]                      d_arburst_0,
    output  [D_AXI_LOCKW-1:0]          d_arlock_0 ,
    output  [3:0]                      d_arcache_0,
    output  [2:0]                      d_arprot_0 ,
    input                              d_arready_0,
    input                              d_rvalid_0 ,
    input   [D_AXI_IDW-1:0]            d_rid_0    ,
    input                              d_rlast_0  ,
    input   [D_AXI_DATA_WID-1:0]       d_rdata_0  ,
    input   [1:0]                      d_rresp_0  ,
    output                             d_rready_0 ,
    output                             d_awvalid_0,
    output  [D_AXI_IDW-1:0]            d_awid_0   ,
    output  [D_AXI_ADDR_WID-1:0]       d_awaddr_0 ,
    output  [D_AXI_LENW-1:0]           d_awlen_0  ,
    output  [2:0]                      d_awsize_0 ,
    output  [1:0]                      d_awburst_0,
    output  [D_AXI_LOCKW-1:0]          d_awlock_0 ,
    output  [3:0]                      d_awcache_0,
    output  [2:0]                      d_awprot_0 ,
    input                              d_awready_0,
    output                             d_wvalid_0 ,
    output                             d_wlast_0  ,
    output  [D_AXI_DATA_WID-1:0]       d_wdata_0  ,
    output  [D_AXI_STRBW-1:0]          d_wstrb_0  ,
    input                              d_wready_0 ,
    input                              d_bvalid_0 ,
    input   [D_AXI_IDW-1:0]            d_bid_0    ,
    input   [1:0]                      d_bresp_0  ,
    output                             d_bready_0 ,

    output                             d_arvalid_1,
    output  [D_AXI_IDW-1:0]            d_arid_1   ,
    output  [D_AXI_ADDR_WID-1:0]       d_araddr_1 ,
    output  [D_AXI_LENW-1:0]           d_arlen_1  ,
    output  [2:0]                      d_arsize_1 ,
    output  [1:0]                      d_arburst_1,
    output  [D_AXI_LOCKW-1:0]          d_arlock_1 ,
    output  [3:0]                      d_arcache_1,
    output  [2:0]                      d_arprot_1 ,
    input                              d_arready_1,
    input                              d_rvalid_1 ,
    input   [D_AXI_IDW-1:0]            d_rid_1    ,
    input                              d_rlast_1  ,
    input   [D_AXI_DATA_WID-1:0]       d_rdata_1  ,
    input   [1:0]                      d_rresp_1  ,
    output                             d_rready_1 ,
    output                             d_awvalid_1,
    output  [D_AXI_IDW-1:0]            d_awid_1   ,
    output  [D_AXI_ADDR_WID-1:0]       d_awaddr_1 ,
    output  [D_AXI_LENW-1:0]           d_awlen_1  ,
    output  [2:0]                      d_awsize_1 ,
    output  [1:0]                      d_awburst_1,
    output  [D_AXI_LOCKW-1:0]          d_awlock_1 ,
    output  [3:0]                      d_awcache_1,
    output  [2:0]                      d_awprot_1 ,
    input                              d_awready_1,
    output                             d_wvalid_1 ,
    output                             d_wlast_1  ,
    output  [D_AXI_DATA_WID-1:0]       d_wdata_1  ,
    output  [D_AXI_STRBW-1:0]          d_wstrb_1  ,
    input                              d_wready_1 ,
    input                              d_bvalid_1 ,
    input   [D_AXI_IDW-1:0]            d_bid_1    ,
    input   [1:0]                      d_bresp_1  ,
    output                             d_bready_1 ,

    //dma axi master interface
    output                                  m_arvalid,
    output [ID_WIDTH-1:0]                   m_arid   ,
    output [AXI_AW-1:0]                     m_araddr ,
    output [AXI_LENW-1:0]                   m_arlen  ,
    output [2:0]                            m_arsize ,
    output [1:0]                            m_arburst,
    output [AXI_LOCKW-1:0]                  m_arlock ,
    output [3:0]                            m_arcache,
    output [2:0]                            m_arprot ,
    input                                   m_arready,
    input                                   m_rvalid ,
    input  [ID_WIDTH-1:0]                   m_rid    ,
    input                                   m_rlast  ,
    input  [AXI_DW-1:0]                     m_rdata  ,
    input  [1:0]                            m_rresp  ,
    output                                  m_rready ,

    input      [11:0]                       cfg_apb_PADDR,
    input      [0:0]                        cfg_apb_PSEL,
    input                                   cfg_apb_PENABLE,
    output                                  cfg_apb_PREADY,
    input                                   cfg_apb_PWRITE,
    input      [3:0]                        cfg_apb_PSTRB,
    input      [2:0]                        cfg_apb_PPROT,
    input      [31:0]                       cfg_apb_PWDATA,
    output     [31:0]                       cfg_apb_PRDATA,
    output                                  cfg_apb_PSLVERR,

    output                                  i_interrupt
);

// AXI slave port
    wire  [ID_WIDTH-1:0]                  s_axi_awid = {ID_WIDTH{1'b0}};
    wire  [AXI_AW-1:0]                    s_axi_awaddr = {AXI_AW{1'b0}};
    wire  [7:0]                           s_axi_awlen = {8{1'b0}};
    wire  [2:0]                           s_axi_awsize = {3{1'b0}};
    wire  [1:0]                           s_axi_awburst = {2{1'b0}};
    wire                                  s_axi_awlock = 1'b0;
    wire  [3:0]                           s_axi_awcache = {4{1'b0}};
    wire  [2:0]                           s_axi_awprot = {3{1'b0}};
    wire                                  s_axi_awvalid = 1'b0;
    wire                                  s_axi_awready;
    wire  [AXI_DW-1:0]                    s_axi_wdata = {AXI_DW{1'b0}};
    wire  [STRB_WIDTH-1:0]                s_axi_wstrb = {STRB_WIDTH{1'b0}};
    wire                                  s_axi_wlast = 1'b0;
    wire                                  s_axi_wvalid = 1'b0;
    wire                                  s_axi_wready;
    wire  [ID_WIDTH-1:0]                  s_axi_bid;
    wire  [1:0]                           s_axi_bresp;
    wire                                  s_axi_bvalid;
    wire                                  s_axi_bready = 1'b1;
    wire  [ID_WIDTH-1:0]                  s_axi_arid = {ID_WIDTH{1'b0}};
    wire  [AXI_AW-1:0]                    s_axi_araddr = {AXI_AW{1'b0}};
    wire  [7:0]                           s_axi_arlen = {8{1'b0}};
    wire  [2:0]                           s_axi_arsize = {3{1'b0}};
    wire  [1:0]                           s_axi_arburst = {2{1'b0}};
    wire                                  s_axi_arlock = 1'b0;
    wire  [3:0]                           s_axi_arcache = {4{1'b0}};
    wire  [2:0]                           s_axi_arprot = {3{1'b0}};
    wire                                  s_axi_arvalid = 1'b0;
    wire                                  s_axi_arready;
    wire  [ID_WIDTH-1:0]                  s_axi_rid;
    wire  [AXI_DW-1:0]                    s_axi_rdata;
    wire  [1:0]                           s_axi_rresp;
    wire                                  s_axi_rlast;
    wire                                  s_axi_rvalid;
    wire                                  s_axi_rready = 1'b1;

recuc U_recuc(
    .clk                                ( clk             ),
    .rst_n                              ( rst_n           ),
    .d_arvalid_0                        ( d_arvalid_0     ),
    .d_arid_0                           ( d_arid_0        ),
    .d_araddr_0                         ( d_araddr_0      ),
    .d_arlen_0                          ( d_arlen_0       ),
    .d_arsize_0                         ( d_arsize_0      ),
    .d_arburst_0                        ( d_arburst_0     ),
    .d_arlock_0                         ( d_arlock_0      ),
    .d_arcache_0                        ( d_arcache_0     ),
    .d_arprot_0                         ( d_arprot_0      ),
    .d_arready_0                        ( d_arready_0     ),
    .d_rvalid_0                         ( d_rvalid_0      ),
    .d_rid_0                            ( d_rid_0         ),
    .d_rlast_0                          ( d_rlast_0       ),
    .d_rdata_0                          ( d_rdata_0       ),
    .d_rresp_0                          ( d_rresp_0       ),
    .d_rready_0                         ( d_rready_0      ),
    .d_awvalid_0                        ( d_awvalid_0     ),
    .d_awid_0                           ( d_awid_0        ),
    .d_awaddr_0                         ( d_awaddr_0      ),
    .d_awlen_0                          ( d_awlen_0       ),
    .d_awsize_0                         ( d_awsize_0      ),
    .d_awburst_0                        ( d_awburst_0     ),
    .d_awlock_0                         ( d_awlock_0      ),
    .d_awcache_0                        ( d_awcache_0     ),
    .d_awprot_0                         ( d_awprot_0      ),
    .d_awready_0                        ( d_awready_0     ),
    .d_wvalid_0                         ( d_wvalid_0      ),
    .d_wlast_0                          ( d_wlast_0       ),
    .d_wdata_0                          ( d_wdata_0       ),
    .d_wstrb_0                          ( d_wstrb_0       ),
    .d_wready_0                         ( d_wready_0      ),
    .d_bvalid_0                         ( d_bvalid_0      ),
    .d_bid_0                            ( d_bid_0         ),
    .d_bresp_0                          ( d_bresp_0       ),
    .d_bready_0                         ( d_bready_0      ),
    .d_arvalid_1                        ( d_arvalid_1     ),
    .d_arid_1                           ( d_arid_1        ),
    .d_araddr_1                         ( d_araddr_1      ),
    .d_arlen_1                          ( d_arlen_1       ),
    .d_arsize_1                         ( d_arsize_1      ),
    .d_arburst_1                        ( d_arburst_1     ),
    .d_arlock_1                         ( d_arlock_1      ),
    .d_arcache_1                        ( d_arcache_1     ),
    .d_arprot_1                         ( d_arprot_1      ),
    .d_arready_1                        ( d_arready_1     ),
    .d_rvalid_1                         ( d_rvalid_1      ),
    .d_rid_1                            ( d_rid_1         ),
    .d_rlast_1                          ( d_rlast_1       ),
    .d_rdata_1                          ( d_rdata_1       ),
    .d_rresp_1                          ( d_rresp_1       ),
    .d_rready_1                         ( d_rready_1      ),
    .d_awvalid_1                        ( d_awvalid_1     ),
    .d_awid_1                           ( d_awid_1        ),
    .d_awaddr_1                         ( d_awaddr_1      ),
    .d_awlen_1                          ( d_awlen_1       ),
    .d_awsize_1                         ( d_awsize_1      ),
    .d_awburst_1                        ( d_awburst_1     ),
    .d_awlock_1                         ( d_awlock_1      ),
    .d_awcache_1                        ( d_awcache_1     ),
    .d_awprot_1                         ( d_awprot_1      ),
    .d_awready_1                        ( d_awready_1     ),
    .d_wvalid_1                         ( d_wvalid_1      ),
    .d_wlast_1                          ( d_wlast_1       ),
    .d_wdata_1                          ( d_wdata_1       ),
    .d_wstrb_1                          ( d_wstrb_1       ),
    .d_wready_1                         ( d_wready_1      ),
    .d_bvalid_1                         ( d_bvalid_1      ),
    .d_bid_1                            ( d_bid_1         ),
    .d_bresp_1                          ( d_bresp_1       ),
    .d_bready_1                         ( d_bready_1      ),
    .s_axi_awid                         ( s_axi_awid      ),
    .s_axi_awaddr                       ( s_axi_awaddr    ),
    .s_axi_awlen                        ( s_axi_awlen     ),
    .s_axi_awsize                       ( s_axi_awsize    ),
    .s_axi_awburst                      ( s_axi_awburst   ),
    .s_axi_awlock                       ( s_axi_awlock    ),
    .s_axi_awcache                      ( s_axi_awcache   ),
    .s_axi_awprot                       ( s_axi_awprot    ),
    .s_axi_awvalid                      ( s_axi_awvalid   ),
    .s_axi_awready                      ( s_axi_awready   ),
    .s_axi_wdata                        ( s_axi_wdata     ),
    .s_axi_wstrb                        ( s_axi_wstrb     ),
    .s_axi_wlast                        ( s_axi_wlast     ),
    .s_axi_wvalid                       ( s_axi_wvalid    ),
    .s_axi_wready                       ( s_axi_wready    ),
    .s_axi_bid                          ( s_axi_bid       ),
    .s_axi_bresp                        ( s_axi_bresp     ),
    .s_axi_bvalid                       ( s_axi_bvalid    ),
    .s_axi_bready                       ( s_axi_bready    ),
    .s_axi_arid                         ( s_axi_arid      ),
    .s_axi_araddr                       ( s_axi_araddr    ),
    .s_axi_arlen                        ( s_axi_arlen     ),
    .s_axi_arsize                       ( s_axi_arsize    ),
    .s_axi_arburst                      ( s_axi_arburst   ),
    .s_axi_arlock                       ( s_axi_arlock    ),
    .s_axi_arcache                      ( s_axi_arcache   ),
    .s_axi_arprot                       ( s_axi_arprot    ),
    .s_axi_arvalid                      ( s_axi_arvalid   ),
    .s_axi_arready                      ( s_axi_arready   ),
    .s_axi_rid                          ( s_axi_rid       ),
    .s_axi_rdata                        ( s_axi_rdata     ),
    .s_axi_rresp                        ( s_axi_rresp     ),
    .s_axi_rlast                        ( s_axi_rlast     ),
    .s_axi_rvalid                       ( s_axi_rvalid    ),
    .s_axi_rready                       ( s_axi_rready    ),
    .m_arvalid                          ( m_arvalid       ),
    .m_arid                             ( m_arid          ),
    .m_araddr                           ( m_araddr        ),
    .m_arlen                            ( m_arlen         ),
    .m_arsize                           ( m_arsize        ),
    .m_arburst                          ( m_arburst       ),
    .m_arlock                           ( m_arlock        ),
    .m_arcache                          ( m_arcache       ),
    .m_arprot                           ( m_arprot        ),
    .m_arready                          ( m_arready       ),
    .m_rvalid                           ( m_rvalid        ),
    .m_rid                              ( m_rid           ),
    .m_rlast                            ( m_rlast         ),
    .m_rdata                            ( m_rdata         ),
    .m_rresp                            ( m_rresp         ),
    .m_rready                           ( m_rready        ),
    .cfg_apb_PADDR                      ( cfg_apb_PADDR   ),
    .cfg_apb_PSEL                       ( cfg_apb_PSEL    ),
    .cfg_apb_PENABLE                    ( cfg_apb_PENABLE ),
    .cfg_apb_PREADY                     ( cfg_apb_PREADY  ),
    .cfg_apb_PWRITE                     ( cfg_apb_PWRITE  ),
    .cfg_apb_PSTRB                      ( cfg_apb_PSTRB   ),
    .cfg_apb_PPROT                      ( cfg_apb_PPROT   ),
    .cfg_apb_PWDATA                     ( cfg_apb_PWDATA  ),
    .cfg_apb_PRDATA                     ( cfg_apb_PRDATA  ),
    .cfg_apb_PSLVERR                    ( cfg_apb_PSLVERR ),
    .i_interrupt                        ( i_interrupt     )
);

endmodule