// 模块功能：数据传输内核模块，用于处理从DMA到NoC的通信。
//          该模块接收配置信号并通过AXI接口和NoC接口进行数据读写操作。
// 数据读写操作：   模块处理来自 AXI 接口的数据读写请求，并通过内部的 FIFO 缓存数据，以匹配处理速度和外部接口的速度。
// 配置与控制：     提供配置接口用于动态设置操作模式，如 FIFO 的阈值设置、outstanding 读写请求的配置等。
// 信号整合与处理：  集成多个控制和数据信号，确保数据一致性和同步。

module idma_data_noc_kernel #(
  parameter DATA_FIFO_DEPTH   = 64    ,
  parameter DATA_FIFO_CNT_WID = 6+1   ,
  parameter ADDR_FIFO_DEPTH   = 32    ,
  parameter ADDR_FIFO_CNT_WID = 5+1   ,

  parameter AXI_DATA_WID      = 256   ,
  parameter AXI_ADDR_WID      = 32    ,
  parameter AXI_IDW           = 4     ,
  parameter AXI_LENW          = 4     ,
  parameter AXI_LOCKW         = 2     ,
  parameter AXI_STRBW         = 32    
)
(
input                              	aclk                    ,
input                              	aresetn                 ,
// =========================== m0 ============================
input    [1:0]                      idma_cfg_ready             ,  // DMA配置就绪信号
//rd channel
input                              	rd_afifo_init              ,  // 读地址FIFO初始化信号 
input                              	rd_dfifo_init              ,  // 读数据FIFO初始化信号
output  [DATA_FIFO_CNT_WID-1: 0]    rd_dfifo_word_cnt          ,  // 读数据FIFO计数
output  [ADDR_FIFO_CNT_WID-1: 0]    rd_afifo_word_cnt          ,  // 读地址FIFO计数
input	[3:0]			                    rd_cfg_outstd              ,  // outstanding 配置
input	     			                    rd_cfg_outstd_en           ,
input                               rd_cfg_cross4k_en          ,  // 读通道跨4K页面使能信号
input                               rd_cfg_arvld_hold_en       ,  // 读通道地址有效保持使能信号
input  [DATA_FIFO_CNT_WID-1:0]      rd_cfg_dfifo_thd           ,  // 读通道的数据FIFO阈值
input                               rd_resi_mode               ,  
input  [AXI_ADDR_WID-1:0]           rd_resi_fmapA_addr         ,
input  [AXI_ADDR_WID-1:0]           rd_resi_fmapB_addr         ,
input  [16-1:0]                     rd_resi_addr_gap           ,
input  [16-1:0]                     rd_resi_loop_num           ,
output  							              rd_done_intr               ,
output  [16-1:0]                    debug_dma_rd_in_cnt        ,
//wr channel
input                              	wr_afifo_init              ,
input                              	wr_dfifo_init              ,
output  [DATA_FIFO_CNT_WID-1: 0]    wr_dfifo_word_cnt          ,
output  [ADDR_FIFO_CNT_WID-1: 0]    wr_afifo_word_cnt          ,
input	  [3:0]			                  wr_cfg_outstd              , 
input	     			                    wr_cfg_outstd_en           ,
input                               wr_cfg_cross4k_en          ,
input                               wr_cfg_arvld_hold_en       ,
input				                        wr_cfg_arvld_hold_olen_en   ,
input  [DATA_FIFO_CNT_WID-1:0]      wr_cfg_dfifo_thd           ,
input                               wr_cfg_strb_force          ,
output  							              wr_done_intr               ,
output [16-1:0]                     debug_dma_wr_out_cnt       ,
//axi interface
output                             	arvalid                  ,
output [AXI_IDW-1:0]               	arid                     ,
output [AXI_ADDR_WID-1:0]           araddr                   ,
output [AXI_LENW-1:0]              	arlen                    ,
output [2:0]                       	arsize                   ,
output [1:0]                       	arburst                  ,
output [AXI_LOCKW-1:0]             	arlock                   ,
output [3:0]                       	arcache                  ,
output [2:0]                       	arprot                   ,
input                              	arready                  ,
input                              	rvalid                   ,
input  [AXI_IDW-1:0]               	rid                      ,
input                              	rlast                    ,
input  [AXI_DATA_WID-1:0]          	rdata                    ,
input  [1:0]                       	rresp                    ,
output                             	rready                   ,
output                             	awvalid                  ,
output [AXI_IDW-1:0]               	awid                     ,
output [AXI_ADDR_WID-1:0]           awaddr                   ,
output [AXI_LENW-1:0]              	awlen                    ,
output [2:0]                       	awsize                   ,
output [1:0]                       	awburst                  ,
output [AXI_LOCKW-1:0]             	awlock                   ,
output [3:0]                       	awcache                  ,
output [2:0]                       	awprot                   ,
input                              	awready                  ,
output                              wvalid                   ,
output  [AXI_IDW-1:0]               wid                      ,
output                              wlast                    ,
output  [AXI_DATA_WID-1:0]          wdata                    ,
output  [AXI_STRBW-1:0]             wstrb                    ,
input                             	wready                   ,
input                               bvalid                   ,
input  [AXI_IDW-1:0]                bid                      ,
input  [1:0]                        bresp                    ,
output                              bready                   ,


// base addr
input  [AXI_ADDR_WID-1:0]           base_addr_0,  //单个32bit，只是对应于一个节点的权重addr
input  [AXI_ADDR_WID-1:0]           base_addr_1,
input  [AXI_ADDR_WID-1:0]           base_addr_2,
input  [AXI_ADDR_WID-1:0]           base_addr_3,
input  [AXI_ADDR_WID-1:0]           base_addr_4,
input  [AXI_ADDR_WID-1:0]           base_addr_5,
input  [AXI_ADDR_WID-1:0]           group_base_addr_0,
input  [AXI_ADDR_WID-1:0]           group_base_addr_1,
input  [AXI_ADDR_WID-1:0]           group_base_addr_2,
input  [AXI_ADDR_WID-1:0]           group_base_addr_3,
input  [AXI_ADDR_WID-1:0]           group_base_addr_4,
input  [AXI_ADDR_WID-1:0]           group_base_addr_5,
input  [AXI_ADDR_WID-1:0]           write_base_addr_0,
input  [AXI_ADDR_WID-1:0]           write_base_addr_1,
input  [AXI_ADDR_WID-1:0]           write_base_addr_2,
input  [AXI_ADDR_WID-1:0]           write_base_addr_3,
input  [AXI_ADDR_WID-1:0]           write_base_addr_4,
input  [AXI_ADDR_WID-1:0]           write_base_addr_5,

// noc ports
output                              data_out_valid   ,
output [AXI_DATA_WID-1:0]           data_out_flit    ,
output                              data_out_last    ,
input                               data_out_ready   ,
input                               data_in_valid    ,
input  [AXI_DATA_WID-1:0]           data_in_flit     ,
input                               data_in_last     ,
output                              data_in_ready    ,
output                              ctrl_out_valid   ,
output [AXI_DATA_WID-1:0]           ctrl_out_flit    ,
output                              ctrl_out_last    ,
input                               ctrl_out_ready   ,
input                               ctrl_in_valid    ,
input  [AXI_DATA_WID-1:0]           ctrl_in_flit     ,
input                               ctrl_in_last     ,
output                              ctrl_in_ready    
);

wire                              	rd_req             ;
wire  [AXI_ADDR_WID-1:0]            rd_addr            ;
wire  [31:0]                     	  rd_num             ;
wire                              	rd_addr_ready      ;
wire                              	rd_data_valid      ;
wire  [AXI_DATA_WID-1:0]            rd_data            ;
wire                              	rd_data_ready      ;
wire  [AXI_STRBW-1:0] 	        	  rd_strb            ;
wire                              	wr_req             ;
wire  [AXI_ADDR_WID-1:0]            wr_addr            ;
wire  [31:0]                     	  wr_num             ;
wire                              	wr_addr_ready      ;
wire                             	  wr_data_valid      ;
wire  [AXI_DATA_WID-1:0]            wr_data            ;
wire                                wr_data_ready      ;
wire  [AXI_STRBW-1:0] 	        	  wr_strb            ;


//处理DMA与NoC之间的数据传输，包括地址、数据流的传递。
idma_data_noc_if#(
    .ADDR_WIDTH     ( AXI_ADDR_WID   ),
    .DATA_WIDTH     ( AXI_DATA_WID   ),
    .STRB_WIDTH     ( AXI_DATA_WID/8 )
)u_idma_data_noc_if(
    .clk            ( aclk           ),
    .rst_n          ( aresetn        ),
    .base_addr_0    ( base_addr_0    ),
    .base_addr_1    ( base_addr_1    ),
    .base_addr_2    ( base_addr_2    ),
    .base_addr_3    ( base_addr_3    ),
    .base_addr_4    ( base_addr_4    ),
    .base_addr_5    ( base_addr_5    ),
    .group_base_addr_0( group_base_addr_0  ),
    .group_base_addr_1( group_base_addr_1  ),
    .group_base_addr_2( group_base_addr_2  ),
    .group_base_addr_3( group_base_addr_3  ),
    .group_base_addr_4( group_base_addr_4  ),
    .group_base_addr_5( group_base_addr_5  ),
    .write_base_addr_0( write_base_addr_0  ),
    .write_base_addr_1( write_base_addr_1  ),
    .write_base_addr_2( write_base_addr_2  ),
    .write_base_addr_3( write_base_addr_3  ),
    .write_base_addr_4( write_base_addr_4  ),
    .write_base_addr_5( write_base_addr_5  ),

    .rd_req            ( rd_req            ),
    .rd_addr           ( rd_addr           ),
    .rd_num            ( rd_num            ),
    .rd_addr_ready     ( rd_addr_ready     ),
    .rd_data_valid     ( rd_data_valid     ),
    .rd_data           ( rd_data           ),
    .rd_data_ready     ( rd_data_ready     ),
    .wr_req            ( wr_req            ),
    .wr_addr           ( wr_addr           ),
    .wr_num            ( wr_num            ),
    .wr_addr_ready     ( wr_addr_ready     ),
    .wr_data_valid     ( wr_data_valid     ),
    .wr_data           ( wr_data           ),
    .wr_data_ready     ( wr_data_ready     ),
    .wr_strb           ( wr_strb           ),
    .wr_done_intr      ( wr_done_intr      ),

    .data_out_valid ( data_out_valid ),
    .data_out_flit  ( data_out_flit  ),
    .data_out_last  ( data_out_last  ),
    .data_out_ready ( data_out_ready ),
    .data_in_valid  ( data_in_valid  ),
    .data_in_flit   ( data_in_flit   ),
    .data_in_last   ( data_in_last   ),
    .data_in_ready  ( data_in_ready  ),
    .ctrl_out_valid ( ctrl_out_valid ),
    .ctrl_out_flit  ( ctrl_out_flit  ),
    .ctrl_out_last  ( ctrl_out_last  ),
    .ctrl_out_ready ( ctrl_out_ready ),
    .ctrl_in_valid  ( ctrl_in_valid  ),
    .ctrl_in_flit   ( ctrl_in_flit   ),
    .ctrl_in_last   ( ctrl_in_last   ),
    .ctrl_in_ready  ( ctrl_in_ready  )
);


// 用于处理DMA与AXI之间的数据同步和传输，处理FIFO的读写操作。
idma_sync_256b_top #(
  .DATA_FIFO_DEPTH        (DATA_FIFO_DEPTH  ),
  .DATA_FIFO_CNT_WID      (DATA_FIFO_CNT_WID),
  .ADDR_FIFO_DEPTH        (ADDR_FIFO_DEPTH  ),
  .ADDR_FIFO_CNT_WID      (ADDR_FIFO_CNT_WID),
  .AXI_DATA_WID           ( AXI_DATA_WID ),
  .AXI_ADDR_WID           ( AXI_ADDR_WID ),
  .AXI_IDW                ( AXI_IDW ),
  .AXI_LENW               ( AXI_LENW ),
  .AXI_LOCKW              ( AXI_LOCKW ),
  .AXI_STRBW              ( AXI_STRBW )
)
u_idma_sync_256b_top(
    .aclk                            ( aclk                               ),
    .aresetn                         ( aresetn                            ),
    .idma_cfg_ready                  ( idma_cfg_ready                     ),
    .rd_afifo_init                   ( rd_afifo_init                      ),
    .rd_dfifo_init                   ( rd_dfifo_init                      ),
    .rd_dfifo_word_cnt               ( rd_dfifo_word_cnt                  ),
    .rd_afifo_word_cnt               ( rd_afifo_word_cnt                  ),
    .rd_cfg_outstd                   ( rd_cfg_outstd                      ),
    .rd_cfg_outstd_en                ( rd_cfg_outstd_en                   ),
    .rd_cfg_cross4k_en               ( rd_cfg_cross4k_en                  ),
    .rd_cfg_arvld_hold_en            ( rd_cfg_arvld_hold_en               ),
    .rd_cfg_dfifo_thd                ( rd_cfg_dfifo_thd                   ),
    .rd_resi_mode                    ( rd_resi_mode                       ),
    .rd_resi_fmapA_addr              ( rd_resi_fmapA_addr                 ),
    .rd_resi_fmapB_addr              ( rd_resi_fmapB_addr                 ),
    .rd_resi_addr_gap                ( rd_resi_addr_gap                   ),
    .rd_resi_loop_num                ( rd_resi_loop_num                   ),
    .wr_afifo_init                   ( wr_afifo_init                      ),
    .wr_dfifo_init                   ( wr_dfifo_init                      ),
    .wr_dfifo_word_cnt               ( wr_dfifo_word_cnt                  ),
    .wr_afifo_word_cnt               ( wr_afifo_word_cnt                  ),
    .wr_cfg_outstd                   ( wr_cfg_outstd                      ),
    .wr_cfg_outstd_en                ( wr_cfg_outstd_en                   ),
    .wr_cfg_cross4k_en               ( wr_cfg_cross4k_en                  ),
    .wr_cfg_arvld_hold_en            ( wr_cfg_arvld_hold_en               ),
    .wr_cfg_arvld_hold_olen_en       ( wr_cfg_arvld_hold_olen_en          ),
    .wr_cfg_dfifo_thd                ( wr_cfg_dfifo_thd                   ),
    .wr_cfg_strb_force               ( wr_cfg_strb_force                  ),
    .rd_req                          ( rd_req                             ),
    .rd_addr                         ( rd_addr                            ),
    .rd_num                          ( rd_num                             ),
    .rd_addr_ready                   ( rd_addr_ready                      ),
    .rd_data_valid                   ( rd_data_valid                      ),
    .rd_data                         ( rd_data                            ),
    .rd_data_ready                   ( rd_data_ready                      ),
    .rd_strb                         ( rd_strb                            ),
    .rd_done_intr                    ( rd_done_intr                       ),
    .debug_dma_rd_in_cnt             ( debug_dma_rd_in_cnt                ),
    .wr_req                          ( wr_req                             ),
    .wr_addr                         ( wr_addr                            ),
    .wr_num                          ( wr_num                             ),
    .wr_addr_ready                   ( wr_addr_ready                      ),
    .wr_data_valid                   ( wr_data_valid                      ),
    .wr_data                         ( wr_data                            ),
    .wr_data_ready                   ( wr_data_ready                      ),
    .wr_strb                         ( wr_strb                            ),
    .wr_done_intr                    ( wr_done_intr                       ),
    .debug_dma_wr_out_cnt            ( debug_dma_wr_out_cnt               ),
    .arvalid                         ( arvalid                            ),
    .arid                            ( arid                               ),
    .araddr                          ( araddr                             ),
    .arlen                           ( arlen                              ),
    .arsize                          ( arsize                             ),
    .arburst                         ( arburst                            ),
    .arlock                          ( arlock                             ),
    .arcache                         ( arcache                            ),
    .arprot                          ( arprot                             ),
    .arready                         ( arready                            ),
    .rvalid                          ( rvalid                             ),
    .rid                             ( rid                                ),
    .rlast                           ( rlast                              ),
    .rdata                           ( rdata                              ),
    .rresp                           ( rresp                              ),
    .rready                          ( rready                             ),
    .awvalid                         ( awvalid                            ),
    .awid                            ( awid                               ),
    .awaddr                          ( awaddr                             ),
    .awlen                           ( awlen                              ),
    .awsize                          ( awsize                             ),
    .awburst                         ( awburst                            ),
    .awlock                          ( awlock                             ),
    .awcache                         ( awcache                            ),
    .awprot                          ( awprot                             ),
    .awready                         ( awready                            ),
    .wvalid                          ( wvalid                             ),
    .wid                             ( wid                                ),
    .wlast                           ( wlast                              ),
    .wdata                           ( wdata                              ),
    .wstrb                           ( wstrb                              ),
    .wready                          ( wready                             ),
    .bvalid                          ( bvalid                             ),
    .bid                             ( bid                                ),
    .bresp                           ( bresp                              ),
    .bready                          ( bready                             )
);

endmodule